LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

ENTITY control IS PORT (

);

ARCHITECTURE arch_ctrl OF control IS BEGIN

END arch_ctrl;