LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;

ENTITY datapath IS PORT (
    
);

ARCHITECTURE arch_dp OF datapath IS BEGIN

END arch_dp;